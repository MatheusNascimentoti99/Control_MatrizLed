// Copyright (C) 1991-2009 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II"
// VERSION		"Version 9.0 Build 132 02/25/2009 SJ Full Version"
// CREATED ON	"Wed Oct 17 09:12:19 2018"

module pbl(
	A,						//ENTRADA 2^0
	B,						//ENTRADA 2^1
	C,						//ENTRADA 2^2
	D,						//ENTRADA 2^3
	clock,					//ENTRADA DO CLOCK DE 32MHz da Placa FPGA 1k 
	COLUA,					//Saida da coluna A
	COLUB,					//Saida da coluna B
	COLUD,					//Saida da coluna D
	COLUE,					//Saida da coluna E
	LIN0,					//Saida da linha 0
	LIN1,					//Saida da linha 1
	LIN2,					//Saida da linha 2
	LIN3,					//Saida da linha 3
	LIN4,					//Saida da linha 4
	LIN5,					//Saida da linha 5
	LIN6,					//Saida da linha 6
	COLUC					//Saida da coluna C
);

//Entradas do circuito
input	A;
input	B;
input	C;
input	D;
input	clock;

//Saidas do circuito
output	COLUA;
output	COLUB;
output	COLUD;
output	COLUE;
output	LIN0;
output	LIN1;
output	LIN2;
output	LIN3;
output	LIN4;
output	LIN5;
output	LIN6;
output	COLUC;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_184;
wire	SYNTHESIZED_WIRE_185;
wire	SYNTHESIZED_WIRE_186;
wire	SYNTHESIZED_WIRE_187;
wire	SYNTHESIZED_WIRE_188;
wire	SYNTHESIZED_WIRE_189;
wire	SYNTHESIZED_WIRE_190;
wire	SYNTHESIZED_WIRE_191;
wire	SYNTHESIZED_WIRE_192;
wire	SYNTHESIZED_WIRE_193;
wire	SYNTHESIZED_WIRE_194;
wire	SYNTHESIZED_WIRE_38;
wire	SYNTHESIZED_WIRE_195;
wire	SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_74;
wire	SYNTHESIZED_WIRE_75;
wire	SYNTHESIZED_WIRE_76;
wire	SYNTHESIZED_WIRE_77;
wire	SYNTHESIZED_WIRE_78;
wire	SYNTHESIZED_WIRE_79;
wire	SYNTHESIZED_WIRE_80;
wire	SYNTHESIZED_WIRE_81;
wire	SYNTHESIZED_WIRE_82;
wire	SYNTHESIZED_WIRE_83;
wire	SYNTHESIZED_WIRE_84;
wire	SYNTHESIZED_WIRE_85;
wire	SYNTHESIZED_WIRE_86;
wire	SYNTHESIZED_WIRE_87;
wire	SYNTHESIZED_WIRE_88;
wire	SYNTHESIZED_WIRE_89;
wire	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_91;
wire	SYNTHESIZED_WIRE_92;
wire	SYNTHESIZED_WIRE_93;
wire	SYNTHESIZED_WIRE_94;
wire	SYNTHESIZED_WIRE_95;
wire	SYNTHESIZED_WIRE_96;
wire	SYNTHESIZED_WIRE_97;
wire	SYNTHESIZED_WIRE_98;
wire	SYNTHESIZED_WIRE_99;
wire	SYNTHESIZED_WIRE_109;
wire	SYNTHESIZED_WIRE_120;
wire	SYNTHESIZED_WIRE_121;
wire	SYNTHESIZED_WIRE_122;
wire	SYNTHESIZED_WIRE_123;
wire	SYNTHESIZED_WIRE_124;
wire	SYNTHESIZED_WIRE_125;
wire	SYNTHESIZED_WIRE_126;
wire	SYNTHESIZED_WIRE_127;
wire	SYNTHESIZED_WIRE_128;
wire	SYNTHESIZED_WIRE_129;
wire	SYNTHESIZED_WIRE_130;
wire	SYNTHESIZED_WIRE_131;
wire	SYNTHESIZED_WIRE_132;
wire	SYNTHESIZED_WIRE_133;
wire	SYNTHESIZED_WIRE_134;
wire	SYNTHESIZED_WIRE_135;
wire	SYNTHESIZED_WIRE_136;
wire	SYNTHESIZED_WIRE_137;
wire	SYNTHESIZED_WIRE_138;
wire	SYNTHESIZED_WIRE_139;
wire	SYNTHESIZED_WIRE_140;
wire	SYNTHESIZED_WIRE_141;
wire	SYNTHESIZED_WIRE_142;
wire	SYNTHESIZED_WIRE_143;
wire	SYNTHESIZED_WIRE_144;
wire	SYNTHESIZED_WIRE_145;
wire	SYNTHESIZED_WIRE_146;
wire	SYNTHESIZED_WIRE_147;
wire	SYNTHESIZED_WIRE_148;
wire	SYNTHESIZED_WIRE_149;
wire	SYNTHESIZED_WIRE_150;
wire	SYNTHESIZED_WIRE_151;
wire	SYNTHESIZED_WIRE_152;
wire	SYNTHESIZED_WIRE_153;
wire	SYNTHESIZED_WIRE_154;
wire	SYNTHESIZED_WIRE_155;
wire	SYNTHESIZED_WIRE_156;
wire	SYNTHESIZED_WIRE_157;
wire	SYNTHESIZED_WIRE_158;
wire	SYNTHESIZED_WIRE_159;
wire	SYNTHESIZED_WIRE_160;
wire	SYNTHESIZED_WIRE_161;
wire	SYNTHESIZED_WIRE_162;
wire	SYNTHESIZED_WIRE_163;
wire	SYNTHESIZED_WIRE_164;
wire	SYNTHESIZED_WIRE_165;
wire	SYNTHESIZED_WIRE_166;
wire	SYNTHESIZED_WIRE_167;
wire	SYNTHESIZED_WIRE_168;
wire	SYNTHESIZED_WIRE_169;
wire	SYNTHESIZED_WIRE_170;
wire	SYNTHESIZED_WIRE_171;
wire	SYNTHESIZED_WIRE_172;
wire	SYNTHESIZED_WIRE_173;
wire	SYNTHESIZED_WIRE_174;
wire	SYNTHESIZED_WIRE_175;
wire	SYNTHESIZED_WIRE_176;
wire	SYNTHESIZED_WIRE_177;
wire	SYNTHESIZED_WIRE_178;
wire	SYNTHESIZED_WIRE_179;
wire	SYNTHESIZED_WIRE_180;
wire	SYNTHESIZED_WIRE_181;
wire	SYNTHESIZED_WIRE_182;
wire	SYNTHESIZED_WIRE_183;

assign	COLUA = SYNTHESIZED_WIRE_190;
assign	COLUB = SYNTHESIZED_WIRE_191;
assign	COLUD = SYNTHESIZED_WIRE_193;
assign	COLUE = SYNTHESIZED_WIRE_194;
assign	COLUC = SYNTHESIZED_WIRE_192;
assign	SYNTHESIZED_WIRE_195 = 1;




Contador3bits	b2v_inst(
	.Clock(SYNTHESIZED_WIRE_0),			//Entrada do clock apos passar pelo divisor de frequencia
	.OUT1(SYNTHESIZED_WIRE_186),		//Valores na saida 2^1, apenas dois valores diferentes
	.OUT2(SYNTHESIZED_WIRE_185),		//Valores na saida 2^2, apenas quatro valores diferentes
	.OUT4(SYNTHESIZED_WIRE_187));		//Valores na saida 2^3, apenas oito valores diferentes


assign	SYNTHESIZED_WIRE_193 = SYNTHESIZED_WIRE_184 & SYNTHESIZED_WIRE_185 & SYNTHESIZED_WIRE_186;

assign	SYNTHESIZED_WIRE_194 = SYNTHESIZED_WIRE_187 & SYNTHESIZED_WIRE_188 & SYNTHESIZED_WIRE_189;

assign	SYNTHESIZED_WIRE_184 =  ~SYNTHESIZED_WIRE_187;

assign	SYNTHESIZED_WIRE_188 =  ~SYNTHESIZED_WIRE_185;

assign	SYNTHESIZED_WIRE_189 =  ~SYNTHESIZED_WIRE_186;

//CI para o caracter 4
char4	b2v_inst15(
	//Seletores
	.A(A),					
	.B(B),
	.C(C),
	.D(D),
	
	//Saidas
	.COL1(SYNTHESIZED_WIRE_190),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.OUT0(SYNTHESIZED_WIRE_84),
	.OUT1(SYNTHESIZED_WIRE_124),
	.OUT2(SYNTHESIZED_WIRE_140),
	.OUT4(SYNTHESIZED_WIRE_156),
	.OUT5(SYNTHESIZED_WIRE_172),
	.OUT6(SYNTHESIZED_WIRE_74));

//CI para o caracter 5
char5	b2v_inst16(
	//Seletores
	.A(A),
	.B(B),
	.C(C),
	.D(D),
	
	//Saidas
	.COL1(SYNTHESIZED_WIRE_190),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.COL5(SYNTHESIZED_WIRE_194),
	.OUT1(SYNTHESIZED_WIRE_125),
	.OUT2(SYNTHESIZED_WIRE_141),
	.OUT4(SYNTHESIZED_WIRE_157),
	.OUT5(SYNTHESIZED_WIRE_173));

//CI para o caracter 7
char7	b2v_inst17(
	.A(A),
	.B(B),
	.C(C),
	.D(D),
	.COL1(SYNTHESIZED_WIRE_190),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.COL5(SYNTHESIZED_WIRE_194),
	.OUT1(SYNTHESIZED_WIRE_128),
	.OUT2(SYNTHESIZED_WIRE_143),
	.OUT3(SYNTHESIZED_WIRE_91),
	.OUT4(SYNTHESIZED_WIRE_159),
	.OUT5(SYNTHESIZED_WIRE_175),
	.OUT6(SYNTHESIZED_WIRE_75));

//CI para o caracter 1
char1	b2v_inst18(
	.A(A),
	.B(B),
	.C(C),
	.D(D),
	.COL1(SYNTHESIZED_WIRE_190),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.OUT0(SYNTHESIZED_WIRE_83),
	.OUT1(SYNTHESIZED_WIRE_121),
	.OUT2(SYNTHESIZED_WIRE_137),
	.OUT3(SYNTHESIZED_WIRE_92),
	.OUT4(SYNTHESIZED_WIRE_153),
	.OUT5(SYNTHESIZED_WIRE_169),
	.OUT6(SYNTHESIZED_WIRE_79));

//CI para o caracter 8
char8	b2v_inst19(
	.A(A),
	.B(B),
	.C(C),
	.D(D),
	.COL1(SYNTHESIZED_WIRE_190),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.COL5(SYNTHESIZED_WIRE_194),
	.OUT0(SYNTHESIZED_WIRE_85),
	.OUT1(SYNTHESIZED_WIRE_129),
	.OUT2(SYNTHESIZED_WIRE_144),
	.OUT3(SYNTHESIZED_WIRE_93),
	.OUT4(SYNTHESIZED_WIRE_160),
	.OUT5(SYNTHESIZED_WIRE_176),
	.OUT6(SYNTHESIZED_WIRE_77));

//CI para o caracter 0
Char0	b2v_inst2(
	.A(A),
	.B(B),
	.C(C),
	.D(D),
	.COL1(SYNTHESIZED_WIRE_190),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.COL5(SYNTHESIZED_WIRE_194),
	.OUT0(SYNTHESIZED_WIRE_82),
	.OUT1(SYNTHESIZED_WIRE_120),
	.OUT2(SYNTHESIZED_WIRE_136),
	.OUT3(SYNTHESIZED_WIRE_90),
	.OUT4(SYNTHESIZED_WIRE_152),
	.OUT5(SYNTHESIZED_WIRE_168),
	.OUT6(SYNTHESIZED_WIRE_76));


freqdiv_0	b2v_inst20(
	.CLK(SYNTHESIZED_WIRE_38),
	
	.G(SYNTHESIZED_WIRE_195),
	
	
	
	.DV16(SYNTHESIZED_WIRE_40));


freqdiv_1	b2v_inst21(
	.CLK(SYNTHESIZED_WIRE_40),
	
	.G(SYNTHESIZED_WIRE_195),
	
	
	
	.DV16(SYNTHESIZED_WIRE_0));

//CI para o caracter 6
char6	b2v_inst22(
	.A(A),
	.B(B),
	.C(C),
	.D(D),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.COL5(SYNTHESIZED_WIRE_194),
	.OUT1(SYNTHESIZED_WIRE_127),
	.OUT2(SYNTHESIZED_WIRE_142),
	.OUT4(SYNTHESIZED_WIRE_158),
	.OUT5(SYNTHESIZED_WIRE_174));

//CI para o caracter 9
char9	b2v_inst23(
	.A(A),
	.B(B),
	.C(C),
	.D(D),
	.COL1(SYNTHESIZED_WIRE_190),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.OUT1(SYNTHESIZED_WIRE_130),
	.OUT2(SYNTHESIZED_WIRE_145),
	.OUT4(SYNTHESIZED_WIRE_161),
	.OUT5(SYNTHESIZED_WIRE_177));

//CI para o caracter A
CharA	b2v_inst24(
	.A(A),
	.B(B),
	.C(C),
	.D(D),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.lin1(SYNTHESIZED_WIRE_126),
	.lin2(SYNTHESIZED_WIRE_146),
	.lin4(SYNTHESIZED_WIRE_162),
	.lin5(SYNTHESIZED_WIRE_178),
	.lin6(SYNTHESIZED_WIRE_78));

//CI para o caracter B
CharB	b2v_inst25(
	.A(A),
	.B(B),
	.C(C),
	.D(D),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.COL5(SYNTHESIZED_WIRE_194),
	.lin0(SYNTHESIZED_WIRE_86),
	.lin1(SYNTHESIZED_WIRE_131),
	.lin2(SYNTHESIZED_WIRE_147),
	.lin3(SYNTHESIZED_WIRE_95),
	.lin4(SYNTHESIZED_WIRE_163),
	.lin5(SYNTHESIZED_WIRE_179),
	.lin6(SYNTHESIZED_WIRE_80));

//CI para o caracter C
CharC	b2v_inst26(
	.A(A),
	.B(B),
	.C(C),
	.D(D),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.COL5(SYNTHESIZED_WIRE_194),
	.lin1(SYNTHESIZED_WIRE_132),
	.lin2(SYNTHESIZED_WIRE_148),
	.lin3(SYNTHESIZED_WIRE_94),
	.lin4(SYNTHESIZED_WIRE_164),
	.lin5(SYNTHESIZED_WIRE_180));

//CI para o caracter D
CharD	b2v_inst27(
	.A(A),
	.B(B),
	.C(C),
	.D(D),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.COL5(SYNTHESIZED_WIRE_194),
	.lin0(SYNTHESIZED_WIRE_87),
	.lin1(SYNTHESIZED_WIRE_133),
	.lin2(SYNTHESIZED_WIRE_149),
	.lin3(SYNTHESIZED_WIRE_96),
	.lin4(SYNTHESIZED_WIRE_165),
	.lin5(SYNTHESIZED_WIRE_181),
	.lin6(SYNTHESIZED_WIRE_81));

//CI para o caracter E
CharE	b2v_inst28(
	.A(A),
	.B(B),
	.C(C),
	.D(D),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.COL5(SYNTHESIZED_WIRE_194),
	.lin1(SYNTHESIZED_WIRE_134),
	.lin2(SYNTHESIZED_WIRE_150),
	.lin3(SYNTHESIZED_WIRE_97),
	.lin4(SYNTHESIZED_WIRE_166),
	.lin5(SYNTHESIZED_WIRE_182));

//CI para o caracter F
CharF	b2v_inst29(
	.A(A),
	.B(B),
	.C(C),
	.D(D),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.COL5(SYNTHESIZED_WIRE_194),
	.lin1(SYNTHESIZED_WIRE_135),
	.lin2(SYNTHESIZED_WIRE_151),
	.liln3(SYNTHESIZED_WIRE_98),
	.lin4(SYNTHESIZED_WIRE_167),
	.lin5(SYNTHESIZED_WIRE_183),
	.lin6(SYNTHESIZED_WIRE_88));


freqdiv_2	b2v_inst3(
	.CLK(clock),
	
	.G(SYNTHESIZED_WIRE_195),
	
	
	
	.DV16(SYNTHESIZED_WIRE_109));

assign	SYNTHESIZED_WIRE_89 = SYNTHESIZED_WIRE_74 | SYNTHESIZED_WIRE_75 | SYNTHESIZED_WIRE_76 | SYNTHESIZED_WIRE_77 | SYNTHESIZED_WIRE_78 | SYNTHESIZED_WIRE_79 | SYNTHESIZED_WIRE_80 | SYNTHESIZED_WIRE_81;

assign	LIN0 = SYNTHESIZED_WIRE_82 | SYNTHESIZED_WIRE_83 | SYNTHESIZED_WIRE_84 | SYNTHESIZED_WIRE_85 | SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_87;

assign	LIN6 = SYNTHESIZED_WIRE_88 | SYNTHESIZED_WIRE_89;

assign	SYNTHESIZED_WIRE_99 = SYNTHESIZED_WIRE_90 | SYNTHESIZED_WIRE_91 | SYNTHESIZED_WIRE_92 | SYNTHESIZED_WIRE_93 | SYNTHESIZED_WIRE_94 | SYNTHESIZED_WIRE_95 | SYNTHESIZED_WIRE_96 | SYNTHESIZED_WIRE_97;

assign	LIN3 = SYNTHESIZED_WIRE_98 | SYNTHESIZED_WIRE_99;

//CI para o caracter 2
char2	b2v_inst4(
	.A(A),
	.B(B),
	.C(C),
	.D(D),
	.COL1(SYNTHESIZED_WIRE_190),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.COL5(SYNTHESIZED_WIRE_194),
	.OUT1(SYNTHESIZED_WIRE_122),
	.OUT2(SYNTHESIZED_WIRE_138),
	.OUT4(SYNTHESIZED_WIRE_154),
	.OUT5(SYNTHESIZED_WIRE_170));

//CI para o caracter 3
char3	b2v_inst5(
	.A(A),
	.B(B),
	.C(C),
	.D(D),
	.COL1(SYNTHESIZED_WIRE_190),
	.COL2(SYNTHESIZED_WIRE_191),
	.COL3(SYNTHESIZED_WIRE_192),
	.COL4(SYNTHESIZED_WIRE_193),
	.OUT1(SYNTHESIZED_WIRE_123),
	.OUT2(SYNTHESIZED_WIRE_139),
	.OUT4(SYNTHESIZED_WIRE_155),
	.OUT5(SYNTHESIZED_WIRE_171));


freqdiv_3	b2v_inst6(
	.CLK(SYNTHESIZED_WIRE_109),
	
	.G(SYNTHESIZED_WIRE_195),
	
	
	
	.DV16(SYNTHESIZED_WIRE_38));

assign	SYNTHESIZED_WIRE_190 = SYNTHESIZED_WIRE_189 & SYNTHESIZED_WIRE_188 & SYNTHESIZED_WIRE_184;

assign	SYNTHESIZED_WIRE_191 = SYNTHESIZED_WIRE_184 & SYNTHESIZED_WIRE_188 & SYNTHESIZED_WIRE_186;

assign	SYNTHESIZED_WIRE_192 = SYNTHESIZED_WIRE_184 & SYNTHESIZED_WIRE_185 & SYNTHESIZED_WIRE_189;


or16	b2v_linha1(
	.input1(SYNTHESIZED_WIRE_120),
	.input2(SYNTHESIZED_WIRE_121),
	.input3(SYNTHESIZED_WIRE_122),
	.input4(SYNTHESIZED_WIRE_123),
	.input5(SYNTHESIZED_WIRE_124),
	.input6(SYNTHESIZED_WIRE_125),
	.input7(SYNTHESIZED_WIRE_126),
	.input8(SYNTHESIZED_WIRE_127),
	.input9(SYNTHESIZED_WIRE_128),
	.input10(SYNTHESIZED_WIRE_129),
	.input11(SYNTHESIZED_WIRE_130),
	.input12(SYNTHESIZED_WIRE_131),
	.input13(SYNTHESIZED_WIRE_132),
	.input14(SYNTHESIZED_WIRE_133),
	.input15(SYNTHESIZED_WIRE_134),
	.input16(SYNTHESIZED_WIRE_135),
	.out(LIN1));


or16	b2v_linha2(
	.input1(SYNTHESIZED_WIRE_136),
	.input2(SYNTHESIZED_WIRE_137),
	.input3(SYNTHESIZED_WIRE_138),
	.input4(SYNTHESIZED_WIRE_139),
	.input5(SYNTHESIZED_WIRE_140),
	.input6(SYNTHESIZED_WIRE_141),
	.input7(SYNTHESIZED_WIRE_142),
	.input8(SYNTHESIZED_WIRE_143),
	.input9(SYNTHESIZED_WIRE_144),
	.input10(SYNTHESIZED_WIRE_145),
	.input11(SYNTHESIZED_WIRE_146),
	.input12(SYNTHESIZED_WIRE_147),
	.input13(SYNTHESIZED_WIRE_148),
	.input14(SYNTHESIZED_WIRE_149),
	.input15(SYNTHESIZED_WIRE_150),
	.input16(SYNTHESIZED_WIRE_151),
	.out(LIN2));


or16	b2v_linha4(
	.input1(SYNTHESIZED_WIRE_152),
	.input2(SYNTHESIZED_WIRE_153),
	.input3(SYNTHESIZED_WIRE_154),
	.input4(SYNTHESIZED_WIRE_155),
	.input5(SYNTHESIZED_WIRE_156),
	.input6(SYNTHESIZED_WIRE_157),
	.input7(SYNTHESIZED_WIRE_158),
	.input8(SYNTHESIZED_WIRE_159),
	.input9(SYNTHESIZED_WIRE_160),
	.input10(SYNTHESIZED_WIRE_161),
	.input11(SYNTHESIZED_WIRE_162),
	.input12(SYNTHESIZED_WIRE_163),
	.input13(SYNTHESIZED_WIRE_164),
	.input14(SYNTHESIZED_WIRE_165),
	.input15(SYNTHESIZED_WIRE_166),
	.input16(SYNTHESIZED_WIRE_167),
	.out(LIN4));


or16	b2v_linha5(
	.input1(SYNTHESIZED_WIRE_168),
	.input2(SYNTHESIZED_WIRE_169),
	.input3(SYNTHESIZED_WIRE_170),
	.input4(SYNTHESIZED_WIRE_171),
	.input5(SYNTHESIZED_WIRE_172),
	.input6(SYNTHESIZED_WIRE_173),
	.input7(SYNTHESIZED_WIRE_174),
	.input8(SYNTHESIZED_WIRE_175),
	.input9(SYNTHESIZED_WIRE_176),
	.input10(SYNTHESIZED_WIRE_177),
	.input11(SYNTHESIZED_WIRE_178),
	.input12(SYNTHESIZED_WIRE_179),
	.input13(SYNTHESIZED_WIRE_180),
	.input14(SYNTHESIZED_WIRE_181),
	.input15(SYNTHESIZED_WIRE_182),
	.input16(SYNTHESIZED_WIRE_183),
	.out(LIN5));


endmodule

module freqdiv_0(CLK,G,DV16);
/* synthesis black_box */

input CLK;
input G;
output DV16;

endmodule

module freqdiv_1(CLK,G,DV16);
/* synthesis black_box */

input CLK;
input G;
output DV16;

endmodule

module freqdiv_2(CLK,G,DV16);
/* synthesis black_box */

input CLK;
input G;
output DV16;

endmodule

module freqdiv_3(CLK,G,DV16);
/* synthesis black_box */

input CLK;
input G;
output DV16;

endmodule
